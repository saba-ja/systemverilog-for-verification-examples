module print_multi_dim_array_tb();

    initial begin
        byte array_2d[4][6]
    end
endmodule